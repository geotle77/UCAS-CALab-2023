`define IDLE    0
`define LOOKUP  1
`define MISS    2
`define REPLACE 3
`define REFILL  4

`define WRBUF_IDLE  0
`define WRBUF_WRITE 1
