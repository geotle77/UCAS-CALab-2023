`ifndef BUS_LEN
    `define BUS_LEN

    `define FS2DS_BUS_LEN 64
    `define DS2ES_BUS_LEN 148
    `define ES2MS_BUS_LEN 71
    `define MS2WS_BUS_LEN 70
    
    `define WB_RF_BUS 38
`endif