`ifndef BUS_LEN
    `define BUS_LEN

    `define FS2DS_BUS_LEN 64
    `define DS2ES_BUS_LEN 156 //
    `define ES2MS_BUS_LEN 90//
    `define MS2WS_BUS_LEN 70
    
    `define ALU_OP_LEN 19
    `define WB_RF_BUS 38
`endif